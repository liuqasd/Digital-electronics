module yxt_2497_7_3(clk_in,rst,auto,Key,clk_out,beep,codeout,low,middle);

input clk_in;   //1MHZ时钟信号
input rst;      //复位信号
input auto;     //自动播放信号
input [13:0]  Key;     //按键信号

output  reg  clk_out;    //分频后输出
output [7:0] codeout;    //数码管信号
output  reg  beep;
output wire [6:0] low;  //表示低音
output wire [6:0] middle;    //表示中音

reg [13:0] tone;           //当前按下的音

yxt_2497_7_1 #(6*3882/2) l1(clk_in,rst,low[0]);
									
yxt_2497_7_1 #(6*3405/2) l2(clk_in,rst,low[1]);
									
yxt_2497_7_1 #(6*3033/2) l3(clk_in,rst,low[2]);
									
yxt_2497_7_1 #(6*2863/2) l4(clk_in,rst,low[3]);
									
yxt_2497_7_1 #(6*2551/2) l5(clk_in,rst,low[4]);
								
yxt_2497_7_1 #(6*2272/2) l6(clk_in,rst,low[5]);
									
yxt_2497_7_1 #(6*2025/2) l7(clk_in,rst,low[6]);
									

yxt_2497_7_1 #(6*1991/2) m1(clk_in,rst,middle[0]);
									
yxt_2497_7_1 #(6*1702/2) m2(clk_in,rst,middle[1]);
									
yxt_2497_7_1 #(6*1516/2) m3(clk_in,rst,middle[2]);
									
yxt_2497_7_1 #(6*1431/2) m4(clk_in,rst,middle[3]);
									
yxt_2497_7_1 #(6*1275/2) m5(clk_in,rst,middle[4]);
									
yxt_2497_7_1 #(6*1136/2) m6(clk_in,rst,middle[5]);
									
yxt_2497_7_1 #(6*1012/2) m7(clk_in,rst,middle[6]);
						  
yxt_2497_7_1 #(6*250000/2)d4(.clk_in(clk_in), .rst(rst), .clk_div(clk_4HZ));//75个音符，需要用7位2进制来表示 
//四分频自动播放音乐

reg [7:0] count;
									
always @(posedge clk_4HZ or negedge rst)  //当自动播放时，count记录最小周期
begin
	if(!rst)
		count   <= 0;
	else
	begin
		if(auto)
		begin
			if(count == 201)
				count <= 0;
			else
				count <= count + 1'b1;
		end
	end
end

always @(posedge clk_in or negedge rst)
begin
	if(!rst)
		tone <= 0;
	else
	begin
		if(!auto)
			begin
				tone <= Key;
			end
			
		else
		begin
		case(count)              //播放歌曲
				 1: tone <= 14'b000_0000_000_0000;// 0
				 2: tone <= 14'b000_0000_000_0000;// 0
				 3: tone <= 14'b000_0000_000_0000;// 0
				 4: tone <= 14'b000_0000_000_0000;// 0
				 5: tone <= 14'b000_0000_000_0000;// 0
				 6: tone <= 14'b000_0000_001_0000;// 1
				 7: tone <= 14'b000_0100_001_0000;// 3
				 8: tone <= 14'b000_0100_000_0100;// 3
				 
				 9: tone <= 14'b000_0000_001_0000;// 3
				10: tone <= 14'b000_0001_000_0000;// 3
				11: tone <= 14'b000_0001_000_0000;// 3
				12: tone <= 14'b000_0001_000_0000;// 3
				13: tone <= 14'b000_0001_000_0000;// 3
				14: tone <= 14'b000_0000_000_0000;// 2
				15: tone <= 14'b000_0000_000_0000;// 1				
				16: tone <= 14'b000_0000_010_0000;// 2
				
				17: tone <= 14'b000_0000_010_0000;// 2
				18: tone <= 14'b000_0001_000_0000;// 3
				19: tone <= 14'b000_0001_000_0000;// 3
				20: tone <= 14'b000_0000_001_0000;// 3
				21: tone <= 14'b000_0000_001_0000;// 0
				22: tone <= 14'b000_0000_001_0000;// 1
	    		23: tone <= 14'b000_0000_001_0000;// 3		
				24: tone <= 14'b000_0000_000_0000;// 3
				
				25: tone <= 14'b000_0000_000_0000;// 3
				26: tone <= 14'b000_0000_010_0000;// 3
				27: tone <= 14'b000_0000_010_0000;// 3
				28: tone <= 14'b000_0000_000_0001;// 3
				29: tone <= 14'b000_0000_000_0010;// 4
				30: tone <= 14'b000_0000_000_0100;// 3
				31: tone <= 14'b000_0000_000_0100;// 5				
				32: tone <= 14'b000_0000_000_0010;// 1
				
				33: tone <= 14'b000_0000_000_0001;// 1
				34: tone <= 14'b000_0000_000_0000;// 1
				35: tone <= 14'b000_0000_000_0010;// 1
				36: tone <= 14'b000_0000_000_0010;// 1
				37: tone <= 14'b000_0000_000_0010;// 0
				38: tone <= 14'b000_0000_000_0010;// 1
				39: tone <= 14'b000_0000_010_0000;// 4
				40: tone <= 14'b000_0000_010_0000;// 4
								
				41: tone <= 14'b000_0000_000_0100;// 4
				42: tone <= 14'b000_0000_001_0000;// 4
				43: tone <= 14'b000_0001_000_0000;// 4
				44: tone <= 14'b000_0001_000_0000;// 4
				45: tone <= 14'b000_0001_000_0000;// 4
				46: tone <= 14'b000_0000_100_0000;// 3
				47: tone <= 14'b000_0000_100_0000;// 1				
				48: tone <= 14'b000_0000_000_0000;//`5
				
				49: tone <= 14'b000_0000_010_0000;//`5
				50: tone <= 14'b000_0000_010_0000;// 3
				51: tone <= 14'b000_0001_000_0000;// 3
				52: tone <= 14'b000_0001_000_0000;// 3
				53: tone <= 14'b000_0000_010_0000;// 0
				54: tone <= 14'b000_0000_010_0000;// 1
				55: tone <= 14'b000_0000_010_0000;// 3
				56: tone <= 14'b000_0000_010_0000;// 2
				
				57: tone <= 14'b000_0000_000_0000;// 2
				58: tone <= 14'b000_0000_000_0000;// 2
				59: tone <= 14'b000_0000_010_0000;// 1
				60: tone <= 14'b000_0000_010_0000;// 3
				61: tone <= 14'b000_0000_000_0010;// 2
				62: tone <= 14'b000_0000_000_0100;// 1
				63: tone <= 14'b000_0000_000_1000;// 3				
				64: tone <= 14'b000_0000_000_1000;// 2
				
				65: tone <= 14'b000_0000_000_1000;// 2
				66: tone <= 14'b000_0000_000_0000;// 2
				67: tone <= 14'b000_0000_000_0001;// 2
				68: tone <= 14'b000_0000_000_0001;// 2
				69: tone <= 14'b000_0000_000_0001;// 0
				70: tone <= 14'b000_0000_000_0001;// 1
//				71: tone <= 14'b000_0100_000_0000;// 3				
//				72: tone <= 14'b000_0100_000_0000;// 3
//				
//				73: tone <= 14'b000_0000_000_0000;// 0
//				74: tone <= 14'b000_0001_000_0000;//`1
//				75: tone <= 14'b000_0001_000_0000;//`1
//				76: tone <= 14'b000_0001_000_0000;//`1
//				77: tone <= 14'b000_0001_000_0000;//`1
//				78: tone <= 14'b000_0000_100_0000;// 7
//				79: tone <= 14'b000_0000_001_0000;// 5				
//				80: tone <= 14'b000_0000_000_0100;// 3
//				
//				81: tone <= 14'b000_0100_000_0000;// 3
//				82: tone <= 14'b000_0100_000_0000;// 3
//				83: tone <= 14'b000_0100_000_0000;// 3 
//				84: tone <= 14'b000_0100_000_0000;// 3
//				85: tone <= 14'b000_0100_000_0000;// 3
//				86: tone <= 14'b000_0010_000_0000;// 2
//				87: tone <= 14'b000_0001_000_0000;// 1				
//				88: tone <= 14'b000_0010_000_0000;// 2
//				
//				89: tone <= 14'b000_0010_000_0000;// 2
//				90: tone <= 14'b001_0000_000_0000;// 5
//				91: tone <= 14'b001_0001_000_0000;// 5
//				92: tone <= 14'b000_0100_000_0000;// 3
//				93: tone <= 14'b000_0000_000_0000;// 0
//				94: tone <= 14'b000_0001_000_0000;// 1
//				95: tone <= 14'b000_0100_000_0000;// 3				
//				96: tone <= 14'b000_0100_000_0000;// 3
//				
//				97: tone <= 14'b000_0100_000_0000;// 3
//				98: tone <= 14'b000_0100_000_0000;// 3
//				99: tone <= 14'b000_0100_000_0000;// 3
//			   100:tone <= 14'b000_0100_000_0000;// 3
//				101:tone <= 14'b000_1000_000_0000;// 4
//				102:tone <= 14'b000_0100_000_0000;// 3
//				103:tone <= 14'b001_0000_000_0000;// 5
//				104:tone <= 14'b000_0001_000_0000;// 1
//				
//				105:tone <= 14'b000_0000_000_0000;// 1
//				106:tone <= 14'b000_0001_000_0000;// 1
//				107:tone <= 14'b000_0001_000_0000;// 1
//				108:tone <= 14'b000_0001_000_0000;// 1
//				109:tone <= 14'b000_0000_000_0000;// 0
//				110:tone <= 14'b000_0001_000_0000;// 1
//				111:tone <= 14'b000_1000_000_0000;// 4
//				112:tone <= 14'b000_1000_000_0000;// 4
//				
//				113:tone <= 14'b000_1000_000_0000;// 4
//				114:tone <= 14'b000_1000_000_0000;// 4
//				115:tone <= 14'b000_1000_000_0000;// 4
//				116:tone <= 14'b000_1000_000_0000;// 4
//				117:tone <= 14'b000_1000_000_0000;// 4
//				118:tone <= 14'b000_0100_000_0000;// 3
//				119:tone <= 14'b000_0001_000_0000;// 1
//				120:tone <= 14'b001_0000_000_0000;// 5
//				
//				121:tone <= 14'b001_0000_000_0000;// 5
//				122:tone <= 14'b000_0100_000_0000;// 3
//				123:tone <= 14'b000_0100_000_0000;// 3
//				124:tone <= 14'b100_0000_000_0000;// 7
//				125:tone <= 14'b100_0000_000_0000;// 7
//				126:tone <= 14'b010_0000_000_0000;// 6
//				127:tone <= 14'b010_0000_000_0000;// 6
//				128:tone <= 14'b000_0000_000_0000;// 0
//				
//				129:tone <= 14'b001_0000_000_0000;// 5
//				130:tone <= 14'b000_1000_000_0000;// 4 
//				131:tone <= 14'b000_1000_000_0000;// 4
//				132:tone <= 14'b000_0001_000_0000;// 1
//				133:tone <= 14'b000_0001_000_0000;// 1
//				134:tone <= 14'b000_0001_000_0000;// 1
//				135:tone <= 14'b000_0000_100_0000;//`7
//				136:tone <= 14'b000_0001_000_0000;// 1
//				
//				137:tone <= 14'b000_0001_000_0000;// 1
//				138:tone <= 14'b000_0001_000_0000;// 1
//				139:tone <= 14'b000_0001_000_0000;// 1
//				140:tone <= 14'b000_0001_000_0000;// 1
//				141:tone <= 14'b000_0010_000_0000;// 2
//				142:tone <= 14'b000_0100_000_0000;// 3
//				143:tone <= 14'b001_0000_000_0000;// 5
//				144:tone <= 14'b001_0000_000_0000;// 5
//				
//				145:tone <= 14'b001_0000_000_0000;// 5
//				146:tone <= 14'b001_0000_000_0000;// 5
//				147:tone <= 14'b001_0000_000_0000;// 5
//				148:tone <= 14'b000_0100_000_0000;// 3
//				149:tone <= 14'b000_0010_000_0000;// 2
//				150:tone <= 14'b000_0001_000_0000;// 1
//				151:tone <= 14'b000_0010_000_0000;// 2
//				152:tone <= 14'b000_0100_000_0000;// 3
//				
//				153:tone <= 14'b000_0100_000_0000;// 3
//				154:tone <= 14'b000_0100_000_0000;// 3
//				155:tone <= 14'b000_0100_000_0000;// 3
//				156:tone <= 14'b000_0100_000_0000;// 3
//				157:tone <= 14'b000_0001_000_0000;// 1
//				158:tone <= 14'b000_0010_000_0000;// 2
//				159:tone <= 14'b000_0100_000_0000;// 3
//				160:tone <= 14'b100_0000_000_0000;// 7
//				
//				161:tone <= 14'b100_0000_000_0000;// 7
//				162:tone <= 14'b100_0000_000_0000;// 7
//				163:tone <= 14'b100_0000_000_0000;// 7
//				164:tone <= 14'b100_0000_000_0000;// 7
//				165:tone <= 14'b010_0000_000_0000;// 6
//				166:tone <= 14'b001_0000_000_0000;// 5
//				167:tone <= 14'b010_0000_000_0000;// 6
//				168:tone <= 14'b010_0000_000_0000;// 6
//				
//				169:tone <= 14'b010_0000_000_0000;// 6
//				170:tone <= 14'b001_0000_000_0000;// 5
//				171:tone <= 14'b001_0000_000_0000;// 5
//				172:tone <= 14'b000_0000_000_0000;// 0
//				173:tone <= 14'b000_0001_000_0000;// 1
//				174:tone <= 14'b000_0010_000_0000;// 2
//				175:tone <= 14'b000_0100_000_0000;// 3
//				176:tone <= 14'b001_0000_000_0000;// 5
//				
//				177:tone <= 14'b001_0000_000_0000;// 5
//				178:tone <= 14'b001_0000_000_0000;// 5
//				179:tone <= 14'b001_0000_000_0000;// 5
//				180:tone <= 14'b000_0100_000_0000;// 3
//				181:tone <= 14'b000_0010_000_0000;// 2
//				182:tone <= 14'b000_0001_000_0000;// 1
//				183:tone <= 14'b000_0010_000_0000;// 2
//				184:tone <= 14'b000_0001_000_0000;// 1
//		
//				185:tone <= 14'b010_0000_000_0000;// 1
//				186:tone <= 14'b001_0000_000_0000;// 1
//				187:tone <= 14'b001_0000_000_0000;// 1
//				188:tone <= 14'b000_0000_000_0000;// 1
//				189:tone <= 14'b000_0001_000_0000;// 1
//				190:tone <= 14'b000_0010_000_0000;// 2
//				191:tone <= 14'b000_0100_000_0000;// 3
//				192:tone <= 14'b001_0000_000_0000;// 5
//
//				193:tone <= 14'b001_0000_000_0000;// 5
//				194:tone <= 14'b000_1000_000_0000;// 4
//				195:tone <= 14'b000_1000_000_0000;// 4
//				196:tone <= 14'b000_0100_000_0000;// 3
//				197:tone <= 14'b100_0000_000_0000;// 7
//				198:tone <= 14'b100_0000_000_0000;// 7
//				199:tone <= 14'b000_0100_000_0000;// 3
//				200:tone <= 14'b000_0100_000_0000;// 3

				71:tone <= 14'b000_0000_000_0001;
				72:tone <= 14'b000_0000_000_0001;
				73:tone <= 14'b000_0000_000_0001;
				74:tone <= 14'b000_0000_000_0001;//7%7+1 = 1
			endcase	
	   end
	end
end


always@(clk_in or tone)      //分频信号始终与当前音对应的频率一致
begin
	case(tone)
		14'b000_0000_000_0000: clk_out <= 0;
		14'b000_0000_000_0001: clk_out <= low[0];
		14'b000_0000_000_0010: clk_out <= low[1];
		14'b000_0000_000_0100: clk_out <= low[2];
		14'b000_0000_000_1000: clk_out <= low[3];
		14'b000_0000_001_0000: clk_out <= low[4];
		14'b000_0000_010_0000: clk_out <= low[5];
		14'b000_0000_100_0000: clk_out <= low[6];
			
		14'b000_0001_000_0000: clk_out <=   middle[0];
		14'b000_0010_000_0000: clk_out <=   middle[1];
		14'b000_0100_000_0000: clk_out <=   middle[2];
		14'b000_1000_000_0000: clk_out <=   middle[3];
		14'b001_0000_000_0000: clk_out <=   middle[4];
		14'b010_0000_000_0000: clk_out <=   middle[5];
		14'b100_0000_000_0000: clk_out <=   middle[6];
	endcase
end
	
always @(clk_in or clk_out)
begin
	beep <= clk_out;
end

yxt_2497_7_2 show(
					   .clk_in(clk_in),
					   .Key(tone),
				   	.codeout(codeout)
				     );
					 
					  
endmodule
