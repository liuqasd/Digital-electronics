module ly_2257_7_3(clk_in,rst,auto,Key,clk_out,clk_out2,codeout,low,middle);

input clk_in;   //时钟信号
input rst;      //复位信号
input auto;     //自动播放信号
input [13:0]  Key;     //按键信号

output reg   clk_out;   //分频后输出
output reg   clk_out2;	//输出频率
output [7:0] codeout;   //数码管信号

output wire  [6:0] low;   	 //表示低音
output wire  [6:0] middle;  //表示中音

reg [13:0] tone;            //当前按下的音

ly_2257_7_1 #(6*3882/2) l1(clk_in,rst,low[0]);
									
ly_2257_7_1 #(6*3405/2) l2(clk_in,rst,low[1]);
									
ly_2257_7_1 #(6*3033/2) l3(clk_in,rst,low[2]);
									
ly_2257_7_1 #(6*2863/2) l4(clk_in,rst,low[3]);
									
ly_2257_7_1 #(6*2551/2) l5(clk_in,rst,low[4]);
								
ly_2257_7_1 #(6*2272/2) l6(clk_in,rst,low[5]);
									
ly_2257_7_1 #(6*2025/2) l7(clk_in,rst,low[6]);
									
									
ly_2257_7_1 #(6*1991/2) m1(clk_in,rst,middle[0]);
									
ly_2257_7_1 #(6*1702/2) m2(clk_in,rst,middle[1]);
									
ly_2257_7_1 #(6*1516/2) m3(clk_in,rst,middle[2]);
									
ly_2257_7_1 #(6*1431/2) m4(clk_in,rst,middle[3]);
									
ly_2257_7_1 #(6*1275/2) m5(clk_in,rst,middle[4]);
									
ly_2257_7_1 #(6*1136/2) m6(clk_in,rst,middle[5]);
									
ly_2257_7_1 #(6*1012/2) m7(clk_in,rst,middle[6]);
						  
ly_2257_7_1 #(6*250000/2)d4(.clk_in(clk_in), .rst(rst), .clk_div(clk_4HZ));//75个音符，需要用7位2进制来表示 
//四分频自动播放音乐

reg [7:0] count;
									
always @(posedge clk_4HZ or negedge rst)  //当自动播放时，count记录最小周期
begin
	if(!rst)
		count   <= 0;
	else
	begin
		if(auto)
		begin
			if(count == 61)	
				count <= 0;
			else
				count <= count + 1'b1;
		end
	end
end

always @(posedge clk_in or negedge rst)
begin
	if(!rst)
		tone <= 0;
	else
	begin
		if(!auto)	tone <= Key;
		else
		begin
			case(count)             //播放《探窗》（C调）
					 1: tone <= 14'b000_0000_000_0000;// 0
					 2: tone <= 14'b000_0100_000_0000;// 3
					 3: tone <= 14'b001_0000_000_0000;// 5
					 4: tone <= 14'b000_0100_000_0000;// 3
					 
					 5: tone <= 14'b000_0010_000_0000;// 2
					 6: tone <= 14'b000_0100_000_0000;// 3
					 7: tone <= 14'b001_0000_000_0000;// 5
					 8: tone <= 14'b000_0100_000_0000;// 3
					 
					 9: tone <= 14'b000_0010_000_0000;// 2
					10: tone <= 14'b000_0010_000_0000;// 2
					11: tone <= 14'b001_0000_000_0000;// 5
					12: tone <= 14'b000_0100_000_0000;// 3
					
					13: tone <= 14'b000_0010_000_0000;// 2
					14: tone <= 14'b000_0100_000_0000;// 3
					15: tone <= 14'b001_0000_000_0000;// 5				
					16: tone <= 14'b000_0010_000_0000;// 2
					
					17: tone <= 14'b000_0001_000_0000;// 1
					18: tone <= 14'b000_0001_000_0000;// 1
					19: tone <= 14'b000_0001_000_0000;// 1
					20: tone <= 14'b000_0010_000_0000;// 2
					
					21: tone <= 14'b000_0100_000_0000;// 3	
					22: tone <= 14'b010_0000_000_0000;// 6
					23: tone <= 14'b010_0000_000_0000;// 6		
					24: tone <= 14'b000_0100_000_0000;// 3
					
					25: tone <= 14'b000_0010_000_0000;// 2
					26: tone <= 14'b000_0010_000_0000;// 2
					27: tone <= 14'b000_0010_000_0000;// 2
					28: tone <= 14'b000_0001_000_0000;// 1
					
					29: tone <= 14'b000_0010_000_0000;// 2
					30: tone <= 14'b000_0100_000_0000;// 3
					31: tone <= 14'b000_0100_000_0000;// 3				
					32: tone <= 14'b001_0000_000_0000;// 5
					
					33: tone <= 14'b000_0100_000_0000;// 3
					34: tone <= 14'b001_0000_000_0000;// 5
					35: tone <= 14'b001_0000_000_0000;// 5
					36: tone <= 14'b000_0100_000_0000;// 3
					
					37: tone <= 14'b000_0010_000_0000;// 2
					38: tone <= 14'b000_0100_000_0000;// 3
					39: tone <= 14'b001_0000_000_0000;// 5
					40: tone <= 14'b000_0100_000_0000;// 3
									
					41: tone <= 14'b000_0010_000_0000;// 2
					42: tone <= 14'b000_0100_000_0000;// 3
					43: tone <= 14'b001_0000_000_0000;// 5
					44: tone <= 14'b000_0100_000_0000;// 3
					
					45: tone <= 14'b000_0000_001_0000;// 5
					46: tone <= 14'b010_0000_000_0000;// 6
					47: tone <= 14'b010_0000_000_0000;// 6		
					48: tone <= 14'b000_0100_000_0000;// 3
					
					49: tone <= 14'b000_0100_000_0000;// 3
					50: tone <= 14'b000_0100_000_0000;// 3
					51: tone <= 14'b000_0010_000_0000;// 2
					52: tone <= 14'b000_0001_000_0000;// 1
					
					53: tone <= 14'b000_0010_000_0000;// 2
					54: tone <= 14'b000_0100_000_0000;// 3
					55: tone <= 14'b000_0010_000_0000;// 2
					56: tone <= 14'b000_0001_000_0000;// 1
					
					
					57: tone <= 14'b000_0010_000_0000;// 2
					58: tone <= 14'b000_0100_000_0000;// 3
					59: tone <= 14'b000_0010_000_0000;// 2
					60: tone <= 14'b010_0000_000_0000;// 6             

					61: tone <= 14'b010_0000_000_0000;// 1 = 7%7+1
			endcase	
	   end
	end
end


always@(clk_in or tone)      //分频信号始终与当前音对应的频率一致
begin
	case(tone)
		14'b000_0000_000_0000: clk_out <= 0;
		14'b000_0000_000_0001: clk_out <= low[0];
		14'b000_0000_000_0010: clk_out <= low[1];
		14'b000_0000_000_0100: clk_out <= low[2];
		14'b000_0000_000_1000: clk_out <= low[3];
		14'b000_0000_001_0000: clk_out <= low[4];
		14'b000_0000_010_0000: clk_out <= low[5];
		14'b000_0000_100_0000: clk_out <= low[6];
			
		14'b000_0001_000_0000: clk_out <= middle[0];
		14'b000_0010_000_0000: clk_out <= middle[1];
		14'b000_0100_000_0000: clk_out <= middle[2];
		14'b000_1000_000_0000: clk_out <= middle[3];
		14'b001_0000_000_0000: clk_out <= middle[4];
		14'b010_0000_000_0000: clk_out <= middle[5];
		14'b100_0000_000_0000: clk_out <= middle[6];
	endcase
end
	
always @(clk_in or clk_out)	clk_out2 <= clk_out;

ly_2257_7_2 show(
	.clk_in(clk_in),
	.Key(tone),
	.codeout(codeout)
);
					 				  
endmodule
